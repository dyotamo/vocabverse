module util

fn test_index() {
	assert true
}
