module util

fn test_web() {
	assert true
}
